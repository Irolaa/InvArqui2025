module Adder8Bit(input [7:0]A,output [7:0]S);
	
logic Ci = 0;
logic [7:0] B = 8'b00000001;	
 logic auxCo1;
 logic auxCo2;
 logic auxCO3;
 logic auxCo4;
 logic auxCo5;
 logic auxCO6;
 logic auxCo7;

 
 
 AdderBit Adder1(A[0], B[0], Ci, auxCo1, S[0]);
 AdderBit Adder2(A[1], B[1], auxCo1, auxCo2, S[1]);
 AdderBit Adder3(A[2], B[2], auxCo2, auxCO3, S[2]);
 AdderBit Adder4(A[3], B[3], auxCO3, auxCo4, S[3]);
 AdderBit Adder5(A[4], B[4], auxCo4, auxCo5, S[4]);
 AdderBit Adder6(A[5], B[5], auxCo5, auxCO6, S[5]);
 AdderBit Adder7(A[6], B[6], auxCO6, auxCo7, S[6]);
 AdderBit Adder8(A[7], B[7], auxCo7, Co, S[7]);

 
 endmodule